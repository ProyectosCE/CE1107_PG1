module Uart_Struct(



);


endmodule 
