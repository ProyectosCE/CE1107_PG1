module FSM_Uart(

);


endmodule 